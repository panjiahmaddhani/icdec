magic
tech sky130A
magscale 1 2
timestamp 1729407255
<< viali >>
rect 3777 2822 3829 2874
rect 3777 2632 3828 2684
rect 3776 2407 3827 2459
<< metal1 >>
rect 3777 2981 3829 2987
rect 900 2920 1247 2955
rect 3777 2923 3829 2929
rect 1212 2865 1247 2920
rect 3765 2874 3841 2880
rect 3765 2865 3777 2874
rect 1212 2831 3777 2865
rect 3119 2678 3153 2831
rect 3765 2822 3777 2831
rect 3829 2822 3841 2874
rect 3765 2816 3841 2822
rect 3766 2727 3776 2779
rect 3828 2727 3838 2779
rect 3771 2684 3834 2696
rect 3771 2675 3777 2684
rect 1210 2624 1503 2659
rect 3614 2641 3777 2675
rect 1106 2130 1158 2136
rect 922 2085 1106 2118
rect 1106 2072 1158 2078
rect 1210 888 1245 2624
rect 3614 1954 3648 2641
rect 3771 2632 3777 2641
rect 3828 2632 3834 2684
rect 3771 2620 3834 2632
rect 3767 2576 3837 2582
rect 3767 2500 3837 2506
rect 3770 2459 3833 2471
rect 3770 2407 3776 2459
rect 3827 2407 3833 2459
rect 3770 2395 3833 2407
rect 3201 1920 3648 1954
rect 1288 1597 1294 1649
rect 1346 1639 1352 1649
rect 1346 1606 1508 1639
rect 1346 1597 1352 1606
rect 2014 1477 2048 1517
rect 1733 1443 2048 1477
rect 1733 1375 1767 1443
rect 901 853 1245 888
rect 2169 268 2203 316
rect 3785 268 3819 2395
rect 2169 234 3819 268
<< via1 >>
rect 3777 2929 3829 2981
rect 3776 2727 3828 2779
rect 1106 2078 1158 2130
rect 3767 2506 3837 2576
rect 1294 1597 1346 1649
<< metal2 >>
rect 2005 2929 3777 2981
rect 3829 2929 3835 2981
rect 2005 2200 2057 2929
rect 3776 2779 3828 2789
rect 3567 2738 3776 2768
rect 1100 2078 1106 2130
rect 1158 2120 1164 2130
rect 1158 2087 1337 2120
rect 3567 2091 3601 2738
rect 3776 2717 3828 2727
rect 1158 2078 1164 2087
rect 1304 1655 1337 2087
rect 3200 2057 3601 2091
rect 3681 2506 3767 2576
rect 3837 2506 3843 2576
rect 3681 1792 3751 2506
rect 3677 1732 3686 1792
rect 3746 1732 3755 1792
rect 3681 1727 3751 1732
rect 1294 1649 1346 1655
rect 1294 1591 1346 1597
rect 2225 1498 2291 1502
rect 892 1493 2296 1498
rect 892 1427 2225 1493
rect 2291 1427 2296 1493
rect 892 1422 2296 1427
rect 2225 1418 2291 1422
rect 2660 1093 2916 1145
rect 2660 880 2712 1093
rect 2375 828 2712 880
<< via2 >>
rect 3686 1732 3746 1792
rect 2225 1427 2291 1493
<< metal3 >>
rect 3681 1792 3751 1797
rect 3681 1732 3686 1792
rect 3746 1732 3751 1792
rect 2220 1493 3176 1498
rect 2220 1427 2225 1493
rect 2291 1427 3176 1493
rect 2220 1422 3176 1427
rect 3681 1153 3751 1732
rect 3356 1093 3751 1153
rect 2367 286 2437 634
rect 3681 286 3751 1093
rect 2367 216 3751 286
use nmos89  nmos89_0
timestamp 1729244476
transform 1 0 1503 0 1 566
box -217 -256 1243 832
use nmoscs  nmoscs_0
timestamp 1729407255
transform 1 0 1630 0 1 1589
box -288 -78 976 1163
use pmos67  pmos67_0
timestamp 1729238107
transform 1 0 2927 0 1 2055
box -197 -1743 621 693
use pmoscs  pmoscs_0
timestamp 1729156831
transform 1 0 249 0 1 833
box -249 -833 916 2158
<< labels >>
flabel via1 3804 2956 3804 2956 0 FreeSans 800 0 0 0 RS
port 0 nsew
flabel viali 3802 2849 3802 2849 0 FreeSans 800 0 0 0 VDD
port 1 nsew
flabel via1 3803 2753 3803 2753 0 FreeSans 800 0 0 0 VIN
port 2 nsew
flabel viali 3802 2659 3802 2659 0 FreeSans 800 0 0 0 VIP
port 3 nsew
flabel via1 3802 2544 3802 2544 0 FreeSans 800 0 0 0 OUT
port 4 nsew
flabel viali 3802 2432 3802 2432 0 FreeSans 800 0 0 0 GND
port 6 nsew
<< end >>
