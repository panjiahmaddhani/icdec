magic
tech sky130A
magscale 1 2
timestamp 1729241244
<< error_p >>
rect -444 345 -372 351
rect -172 345 -100 351
rect 100 345 172 351
rect 372 345 444 351
rect -444 311 -432 345
rect -172 311 -160 345
rect 100 311 112 345
rect 372 311 384 345
rect -444 305 -372 311
rect -172 305 -100 311
rect 100 305 172 311
rect 372 305 444 311
rect -444 17 -372 23
rect -172 17 -100 23
rect 100 17 172 23
rect 372 17 444 23
rect -444 -17 -432 17
rect -172 -17 -160 17
rect 100 -17 112 17
rect 372 -17 384 17
rect -444 -23 -372 -17
rect -172 -23 -100 -17
rect 100 -23 172 -17
rect 372 -23 444 -17
rect -444 -311 -372 -305
rect -172 -311 -100 -305
rect 100 -311 172 -305
rect 372 -311 444 -305
rect -444 -345 -432 -311
rect -172 -345 -160 -311
rect 100 -345 112 -311
rect 372 -345 384 -311
rect -444 -351 -372 -345
rect -172 -351 -100 -345
rect 100 -351 172 -345
rect 372 -351 444 -345
<< nwell >>
rect -552 -364 552 364
<< pmos >>
rect -458 64 -358 264
rect -186 64 -86 264
rect 86 64 186 264
rect 358 64 458 264
rect -458 -264 -358 -64
rect -186 -264 -86 -64
rect 86 -264 186 -64
rect 358 -264 458 -64
<< pdiff >>
rect -516 252 -458 264
rect -516 76 -504 252
rect -470 76 -458 252
rect -516 64 -458 76
rect -358 252 -300 264
rect -358 76 -346 252
rect -312 76 -300 252
rect -358 64 -300 76
rect -244 252 -186 264
rect -244 76 -232 252
rect -198 76 -186 252
rect -244 64 -186 76
rect -86 252 -28 264
rect -86 76 -74 252
rect -40 76 -28 252
rect -86 64 -28 76
rect 28 252 86 264
rect 28 76 40 252
rect 74 76 86 252
rect 28 64 86 76
rect 186 252 244 264
rect 186 76 198 252
rect 232 76 244 252
rect 186 64 244 76
rect 300 252 358 264
rect 300 76 312 252
rect 346 76 358 252
rect 300 64 358 76
rect 458 252 516 264
rect 458 76 470 252
rect 504 76 516 252
rect 458 64 516 76
rect -516 -76 -458 -64
rect -516 -252 -504 -76
rect -470 -252 -458 -76
rect -516 -264 -458 -252
rect -358 -76 -300 -64
rect -358 -252 -346 -76
rect -312 -252 -300 -76
rect -358 -264 -300 -252
rect -244 -76 -186 -64
rect -244 -252 -232 -76
rect -198 -252 -186 -76
rect -244 -264 -186 -252
rect -86 -76 -28 -64
rect -86 -252 -74 -76
rect -40 -252 -28 -76
rect -86 -264 -28 -252
rect 28 -76 86 -64
rect 28 -252 40 -76
rect 74 -252 86 -76
rect 28 -264 86 -252
rect 186 -76 244 -64
rect 186 -252 198 -76
rect 232 -252 244 -76
rect 186 -264 244 -252
rect 300 -76 358 -64
rect 300 -252 312 -76
rect 346 -252 358 -76
rect 300 -264 358 -252
rect 458 -76 516 -64
rect 458 -252 470 -76
rect 504 -252 516 -76
rect 458 -264 516 -252
<< pdiffc >>
rect -504 76 -470 252
rect -346 76 -312 252
rect -232 76 -198 252
rect -74 76 -40 252
rect 40 76 74 252
rect 198 76 232 252
rect 312 76 346 252
rect 470 76 504 252
rect -504 -252 -470 -76
rect -346 -252 -312 -76
rect -232 -252 -198 -76
rect -74 -252 -40 -76
rect 40 -252 74 -76
rect 198 -252 232 -76
rect 312 -252 346 -76
rect 470 -252 504 -76
<< poly >>
rect -458 345 -358 361
rect -458 311 -442 345
rect -374 311 -358 345
rect -458 264 -358 311
rect -186 345 -86 361
rect -186 311 -170 345
rect -102 311 -86 345
rect -186 264 -86 311
rect 86 345 186 361
rect 86 311 102 345
rect 170 311 186 345
rect 86 264 186 311
rect 358 345 458 361
rect 358 311 374 345
rect 442 311 458 345
rect 358 264 458 311
rect -458 17 -358 64
rect -458 -17 -442 17
rect -374 -17 -358 17
rect -458 -64 -358 -17
rect -186 17 -86 64
rect -186 -17 -170 17
rect -102 -17 -86 17
rect -186 -64 -86 -17
rect 86 17 186 64
rect 86 -17 102 17
rect 170 -17 186 17
rect 86 -64 186 -17
rect 358 17 458 64
rect 358 -17 374 17
rect 442 -17 458 17
rect 358 -64 458 -17
rect -458 -311 -358 -264
rect -458 -345 -442 -311
rect -374 -345 -358 -311
rect -458 -361 -358 -345
rect -186 -311 -86 -264
rect -186 -345 -170 -311
rect -102 -345 -86 -311
rect -186 -361 -86 -345
rect 86 -311 186 -264
rect 86 -345 102 -311
rect 170 -345 186 -311
rect 86 -361 186 -345
rect 358 -311 458 -264
rect 358 -345 374 -311
rect 442 -345 458 -311
rect 358 -361 458 -345
<< polycont >>
rect -442 311 -374 345
rect -170 311 -102 345
rect 102 311 170 345
rect 374 311 442 345
rect -442 -17 -374 17
rect -170 -17 -102 17
rect 102 -17 170 17
rect 374 -17 442 17
rect -442 -345 -374 -311
rect -170 -345 -102 -311
rect 102 -345 170 -311
rect 374 -345 442 -311
<< locali >>
rect -458 311 -442 345
rect -374 311 -358 345
rect -186 311 -170 345
rect -102 311 -86 345
rect 86 311 102 345
rect 170 311 186 345
rect 358 311 374 345
rect 442 311 458 345
rect -504 252 -470 268
rect -504 60 -470 76
rect -346 252 -312 268
rect -346 60 -312 76
rect -232 252 -198 268
rect -232 60 -198 76
rect -74 252 -40 268
rect -74 60 -40 76
rect 40 252 74 268
rect 40 60 74 76
rect 198 252 232 268
rect 198 60 232 76
rect 312 252 346 268
rect 312 60 346 76
rect 470 252 504 268
rect 470 60 504 76
rect -458 -17 -442 17
rect -374 -17 -358 17
rect -186 -17 -170 17
rect -102 -17 -86 17
rect 86 -17 102 17
rect 170 -17 186 17
rect 358 -17 374 17
rect 442 -17 458 17
rect -504 -76 -470 -60
rect -504 -268 -470 -252
rect -346 -76 -312 -60
rect -346 -268 -312 -252
rect -232 -76 -198 -60
rect -232 -268 -198 -252
rect -74 -76 -40 -60
rect -74 -268 -40 -252
rect 40 -76 74 -60
rect 40 -268 74 -252
rect 198 -76 232 -60
rect 198 -268 232 -252
rect 312 -76 346 -60
rect 312 -268 346 -252
rect 470 -76 504 -60
rect 470 -268 504 -252
rect -458 -345 -442 -311
rect -374 -345 -358 -311
rect -186 -345 -170 -311
rect -102 -345 -86 -311
rect 86 -345 102 -311
rect 170 -345 186 -311
rect 358 -345 374 -311
rect 442 -345 458 -311
<< viali >>
rect -432 311 -384 345
rect -160 311 -112 345
rect 112 311 160 345
rect 384 311 432 345
rect -504 76 -470 252
rect -346 76 -312 252
rect -232 76 -198 252
rect -74 76 -40 252
rect 40 76 74 252
rect 198 76 232 252
rect 312 76 346 252
rect 470 76 504 252
rect -432 -17 -384 17
rect -160 -17 -112 17
rect 112 -17 160 17
rect 384 -17 432 17
rect -504 -252 -470 -76
rect -346 -252 -312 -76
rect -232 -252 -198 -76
rect -74 -252 -40 -76
rect 40 -252 74 -76
rect 198 -252 232 -76
rect 312 -252 346 -76
rect 470 -252 504 -76
rect -432 -345 -384 -311
rect -160 -345 -112 -311
rect 112 -345 160 -311
rect 384 -345 432 -311
<< metal1 >>
rect -444 345 -372 351
rect -444 311 -432 345
rect -384 311 -372 345
rect -444 305 -372 311
rect -172 345 -100 351
rect -172 311 -160 345
rect -112 311 -100 345
rect -172 305 -100 311
rect 100 345 172 351
rect 100 311 112 345
rect 160 311 172 345
rect 100 305 172 311
rect 372 345 444 351
rect 372 311 384 345
rect 432 311 444 345
rect 372 305 444 311
rect -510 252 -464 264
rect -510 76 -504 252
rect -470 76 -464 252
rect -510 64 -464 76
rect -352 252 -306 264
rect -352 76 -346 252
rect -312 76 -306 252
rect -352 64 -306 76
rect -238 252 -192 264
rect -238 76 -232 252
rect -198 76 -192 252
rect -238 64 -192 76
rect -80 252 -34 264
rect -80 76 -74 252
rect -40 76 -34 252
rect -80 64 -34 76
rect 34 252 80 264
rect 34 76 40 252
rect 74 76 80 252
rect 34 64 80 76
rect 192 252 238 264
rect 192 76 198 252
rect 232 76 238 252
rect 192 64 238 76
rect 306 252 352 264
rect 306 76 312 252
rect 346 76 352 252
rect 306 64 352 76
rect 464 252 510 264
rect 464 76 470 252
rect 504 76 510 252
rect 464 64 510 76
rect -444 17 -372 23
rect -444 -17 -432 17
rect -384 -17 -372 17
rect -444 -23 -372 -17
rect -172 17 -100 23
rect -172 -17 -160 17
rect -112 -17 -100 17
rect -172 -23 -100 -17
rect 100 17 172 23
rect 100 -17 112 17
rect 160 -17 172 17
rect 100 -23 172 -17
rect 372 17 444 23
rect 372 -17 384 17
rect 432 -17 444 17
rect 372 -23 444 -17
rect -510 -76 -464 -64
rect -510 -252 -504 -76
rect -470 -252 -464 -76
rect -510 -264 -464 -252
rect -352 -76 -306 -64
rect -352 -252 -346 -76
rect -312 -252 -306 -76
rect -352 -264 -306 -252
rect -238 -76 -192 -64
rect -238 -252 -232 -76
rect -198 -252 -192 -76
rect -238 -264 -192 -252
rect -80 -76 -34 -64
rect -80 -252 -74 -76
rect -40 -252 -34 -76
rect -80 -264 -34 -252
rect 34 -76 80 -64
rect 34 -252 40 -76
rect 74 -252 80 -76
rect 34 -264 80 -252
rect 192 -76 238 -64
rect 192 -252 198 -76
rect 232 -252 238 -76
rect 192 -264 238 -252
rect 306 -76 352 -64
rect 306 -252 312 -76
rect 346 -252 352 -76
rect 306 -264 352 -252
rect 464 -76 510 -64
rect 464 -252 470 -76
rect 504 -252 510 -76
rect 464 -264 510 -252
rect -444 -311 -372 -305
rect -444 -345 -432 -311
rect -384 -345 -372 -311
rect -444 -351 -372 -345
rect -172 -311 -100 -305
rect -172 -345 -160 -311
rect -112 -345 -100 -311
rect -172 -351 -100 -345
rect 100 -311 172 -305
rect 100 -345 112 -311
rect 160 -345 172 -311
rect 100 -351 172 -345
rect 372 -311 444 -305
rect 372 -345 384 -311
rect 432 -345 444 -311
rect 372 -351 444 -345
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.5 m 2 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 70 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
