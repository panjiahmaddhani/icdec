magic
tech sky130A
magscale 1 2
timestamp 1729241244
<< error_p >>
rect -273 345 -201 351
rect -115 345 -43 351
rect 43 345 115 351
rect 201 345 273 351
rect -273 311 -261 345
rect -115 311 -103 345
rect 43 311 55 345
rect 201 311 213 345
rect -273 305 -201 311
rect -115 305 -43 311
rect 43 305 115 311
rect 201 305 273 311
rect -273 17 -201 23
rect -115 17 -43 23
rect 43 17 115 23
rect 201 17 273 23
rect -273 -17 -261 17
rect -115 -17 -103 17
rect 43 -17 55 17
rect 201 -17 213 17
rect -273 -23 -201 -17
rect -115 -23 -43 -17
rect 43 -23 115 -17
rect 201 -23 273 -17
rect -273 -311 -201 -305
rect -115 -311 -43 -305
rect 43 -311 115 -305
rect 201 -311 273 -305
rect -273 -345 -261 -311
rect -115 -345 -103 -311
rect 43 -345 55 -311
rect 201 -345 213 -311
rect -273 -351 -201 -345
rect -115 -351 -43 -345
rect 43 -351 115 -345
rect 201 -351 273 -345
<< nwell >>
rect -381 -364 381 364
<< pmos >>
rect -287 64 -187 264
rect -129 64 -29 264
rect 29 64 129 264
rect 187 64 287 264
rect -287 -264 -187 -64
rect -129 -264 -29 -64
rect 29 -264 129 -64
rect 187 -264 287 -64
<< pdiff >>
rect -345 252 -287 264
rect -345 76 -333 252
rect -299 76 -287 252
rect -345 64 -287 76
rect -187 252 -129 264
rect -187 76 -175 252
rect -141 76 -129 252
rect -187 64 -129 76
rect -29 252 29 264
rect -29 76 -17 252
rect 17 76 29 252
rect -29 64 29 76
rect 129 252 187 264
rect 129 76 141 252
rect 175 76 187 252
rect 129 64 187 76
rect 287 252 345 264
rect 287 76 299 252
rect 333 76 345 252
rect 287 64 345 76
rect -345 -76 -287 -64
rect -345 -252 -333 -76
rect -299 -252 -287 -76
rect -345 -264 -287 -252
rect -187 -76 -129 -64
rect -187 -252 -175 -76
rect -141 -252 -129 -76
rect -187 -264 -129 -252
rect -29 -76 29 -64
rect -29 -252 -17 -76
rect 17 -252 29 -76
rect -29 -264 29 -252
rect 129 -76 187 -64
rect 129 -252 141 -76
rect 175 -252 187 -76
rect 129 -264 187 -252
rect 287 -76 345 -64
rect 287 -252 299 -76
rect 333 -252 345 -76
rect 287 -264 345 -252
<< pdiffc >>
rect -333 76 -299 252
rect -175 76 -141 252
rect -17 76 17 252
rect 141 76 175 252
rect 299 76 333 252
rect -333 -252 -299 -76
rect -175 -252 -141 -76
rect -17 -252 17 -76
rect 141 -252 175 -76
rect 299 -252 333 -76
<< poly >>
rect -287 345 -187 361
rect -287 311 -271 345
rect -203 311 -187 345
rect -287 264 -187 311
rect -129 345 -29 361
rect -129 311 -113 345
rect -45 311 -29 345
rect -129 264 -29 311
rect 29 345 129 361
rect 29 311 45 345
rect 113 311 129 345
rect 29 264 129 311
rect 187 345 287 361
rect 187 311 203 345
rect 271 311 287 345
rect 187 264 287 311
rect -287 17 -187 64
rect -287 -17 -271 17
rect -203 -17 -187 17
rect -287 -64 -187 -17
rect -129 17 -29 64
rect -129 -17 -113 17
rect -45 -17 -29 17
rect -129 -64 -29 -17
rect 29 17 129 64
rect 29 -17 45 17
rect 113 -17 129 17
rect 29 -64 129 -17
rect 187 17 287 64
rect 187 -17 203 17
rect 271 -17 287 17
rect 187 -64 287 -17
rect -287 -311 -187 -264
rect -287 -345 -271 -311
rect -203 -345 -187 -311
rect -287 -361 -187 -345
rect -129 -311 -29 -264
rect -129 -345 -113 -311
rect -45 -345 -29 -311
rect -129 -361 -29 -345
rect 29 -311 129 -264
rect 29 -345 45 -311
rect 113 -345 129 -311
rect 29 -361 129 -345
rect 187 -311 287 -264
rect 187 -345 203 -311
rect 271 -345 287 -311
rect 187 -361 287 -345
<< polycont >>
rect -271 311 -203 345
rect -113 311 -45 345
rect 45 311 113 345
rect 203 311 271 345
rect -271 -17 -203 17
rect -113 -17 -45 17
rect 45 -17 113 17
rect 203 -17 271 17
rect -271 -345 -203 -311
rect -113 -345 -45 -311
rect 45 -345 113 -311
rect 203 -345 271 -311
<< locali >>
rect -287 311 -271 345
rect -203 311 -187 345
rect -129 311 -113 345
rect -45 311 -29 345
rect 29 311 45 345
rect 113 311 129 345
rect 187 311 203 345
rect 271 311 287 345
rect -333 252 -299 268
rect -333 60 -299 76
rect -175 252 -141 268
rect -175 60 -141 76
rect -17 252 17 268
rect -17 60 17 76
rect 141 252 175 268
rect 141 60 175 76
rect 299 252 333 268
rect 299 60 333 76
rect -287 -17 -271 17
rect -203 -17 -187 17
rect -129 -17 -113 17
rect -45 -17 -29 17
rect 29 -17 45 17
rect 113 -17 129 17
rect 187 -17 203 17
rect 271 -17 287 17
rect -333 -76 -299 -60
rect -333 -268 -299 -252
rect -175 -76 -141 -60
rect -175 -268 -141 -252
rect -17 -76 17 -60
rect -17 -268 17 -252
rect 141 -76 175 -60
rect 141 -268 175 -252
rect 299 -76 333 -60
rect 299 -268 333 -252
rect -287 -345 -271 -311
rect -203 -345 -187 -311
rect -129 -345 -113 -311
rect -45 -345 -29 -311
rect 29 -345 45 -311
rect 113 -345 129 -311
rect 187 -345 203 -311
rect 271 -345 287 -311
<< viali >>
rect -261 311 -213 345
rect -103 311 -55 345
rect 55 311 103 345
rect 213 311 261 345
rect -333 76 -299 252
rect -175 76 -141 252
rect -17 76 17 252
rect 141 76 175 252
rect 299 76 333 252
rect -261 -17 -213 17
rect -103 -17 -55 17
rect 55 -17 103 17
rect 213 -17 261 17
rect -333 -252 -299 -76
rect -175 -252 -141 -76
rect -17 -252 17 -76
rect 141 -252 175 -76
rect 299 -252 333 -76
rect -261 -345 -213 -311
rect -103 -345 -55 -311
rect 55 -345 103 -311
rect 213 -345 261 -311
<< metal1 >>
rect -273 345 -201 351
rect -273 311 -261 345
rect -213 311 -201 345
rect -273 305 -201 311
rect -115 345 -43 351
rect -115 311 -103 345
rect -55 311 -43 345
rect -115 305 -43 311
rect 43 345 115 351
rect 43 311 55 345
rect 103 311 115 345
rect 43 305 115 311
rect 201 345 273 351
rect 201 311 213 345
rect 261 311 273 345
rect 201 305 273 311
rect -339 252 -293 264
rect -339 76 -333 252
rect -299 76 -293 252
rect -339 64 -293 76
rect -181 252 -135 264
rect -181 76 -175 252
rect -141 76 -135 252
rect -181 64 -135 76
rect -23 252 23 264
rect -23 76 -17 252
rect 17 76 23 252
rect -23 64 23 76
rect 135 252 181 264
rect 135 76 141 252
rect 175 76 181 252
rect 135 64 181 76
rect 293 252 339 264
rect 293 76 299 252
rect 333 76 339 252
rect 293 64 339 76
rect -273 17 -201 23
rect -273 -17 -261 17
rect -213 -17 -201 17
rect -273 -23 -201 -17
rect -115 17 -43 23
rect -115 -17 -103 17
rect -55 -17 -43 17
rect -115 -23 -43 -17
rect 43 17 115 23
rect 43 -17 55 17
rect 103 -17 115 17
rect 43 -23 115 -17
rect 201 17 273 23
rect 201 -17 213 17
rect 261 -17 273 17
rect 201 -23 273 -17
rect -339 -76 -293 -64
rect -339 -252 -333 -76
rect -299 -252 -293 -76
rect -339 -264 -293 -252
rect -181 -76 -135 -64
rect -181 -252 -175 -76
rect -141 -252 -135 -76
rect -181 -264 -135 -252
rect -23 -76 23 -64
rect -23 -252 -17 -76
rect 17 -252 23 -76
rect -23 -264 23 -252
rect 135 -76 181 -64
rect 135 -252 141 -76
rect 175 -252 181 -76
rect 135 -264 181 -252
rect 293 -76 339 -64
rect 293 -252 299 -76
rect 333 -252 339 -76
rect 293 -264 339 -252
rect -273 -311 -201 -305
rect -273 -345 -261 -311
rect -213 -345 -201 -311
rect -273 -351 -201 -345
rect -115 -311 -43 -305
rect -115 -345 -103 -311
rect -55 -345 -43 -311
rect -115 -351 -43 -345
rect 43 -311 115 -305
rect 43 -345 55 -311
rect 103 -345 115 -311
rect 43 -351 115 -345
rect 201 -311 273 -305
rect 201 -345 213 -311
rect 261 -345 273 -311
rect 201 -351 273 -345
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.5 m 2 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 70 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
