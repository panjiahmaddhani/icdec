magic
tech sky130A
magscale 1 2
timestamp 1729241244
<< error_p >>
rect -172 673 -100 679
rect 100 673 172 679
rect -172 639 -160 673
rect 100 639 112 673
rect -172 633 -100 639
rect 100 633 172 639
rect -172 345 -100 351
rect 100 345 172 351
rect -172 311 -160 345
rect 100 311 112 345
rect -172 305 -100 311
rect 100 305 172 311
rect -172 17 -100 23
rect 100 17 172 23
rect -172 -17 -160 17
rect 100 -17 112 17
rect -172 -23 -100 -17
rect 100 -23 172 -17
rect -172 -311 -100 -305
rect 100 -311 172 -305
rect -172 -345 -160 -311
rect 100 -345 112 -311
rect -172 -351 -100 -345
rect 100 -351 172 -345
rect -172 -639 -100 -633
rect 100 -639 172 -633
rect -172 -673 -160 -639
rect 100 -673 112 -639
rect -172 -679 -100 -673
rect 100 -679 172 -673
<< nwell >>
rect -280 -692 280 692
<< pmos >>
rect -186 392 -86 592
rect 86 392 186 592
rect -186 64 -86 264
rect 86 64 186 264
rect -186 -264 -86 -64
rect 86 -264 186 -64
rect -186 -592 -86 -392
rect 86 -592 186 -392
<< pdiff >>
rect -244 580 -186 592
rect -244 404 -232 580
rect -198 404 -186 580
rect -244 392 -186 404
rect -86 580 -28 592
rect -86 404 -74 580
rect -40 404 -28 580
rect -86 392 -28 404
rect 28 580 86 592
rect 28 404 40 580
rect 74 404 86 580
rect 28 392 86 404
rect 186 580 244 592
rect 186 404 198 580
rect 232 404 244 580
rect 186 392 244 404
rect -244 252 -186 264
rect -244 76 -232 252
rect -198 76 -186 252
rect -244 64 -186 76
rect -86 252 -28 264
rect -86 76 -74 252
rect -40 76 -28 252
rect -86 64 -28 76
rect 28 252 86 264
rect 28 76 40 252
rect 74 76 86 252
rect 28 64 86 76
rect 186 252 244 264
rect 186 76 198 252
rect 232 76 244 252
rect 186 64 244 76
rect -244 -76 -186 -64
rect -244 -252 -232 -76
rect -198 -252 -186 -76
rect -244 -264 -186 -252
rect -86 -76 -28 -64
rect -86 -252 -74 -76
rect -40 -252 -28 -76
rect -86 -264 -28 -252
rect 28 -76 86 -64
rect 28 -252 40 -76
rect 74 -252 86 -76
rect 28 -264 86 -252
rect 186 -76 244 -64
rect 186 -252 198 -76
rect 232 -252 244 -76
rect 186 -264 244 -252
rect -244 -404 -186 -392
rect -244 -580 -232 -404
rect -198 -580 -186 -404
rect -244 -592 -186 -580
rect -86 -404 -28 -392
rect -86 -580 -74 -404
rect -40 -580 -28 -404
rect -86 -592 -28 -580
rect 28 -404 86 -392
rect 28 -580 40 -404
rect 74 -580 86 -404
rect 28 -592 86 -580
rect 186 -404 244 -392
rect 186 -580 198 -404
rect 232 -580 244 -404
rect 186 -592 244 -580
<< pdiffc >>
rect -232 404 -198 580
rect -74 404 -40 580
rect 40 404 74 580
rect 198 404 232 580
rect -232 76 -198 252
rect -74 76 -40 252
rect 40 76 74 252
rect 198 76 232 252
rect -232 -252 -198 -76
rect -74 -252 -40 -76
rect 40 -252 74 -76
rect 198 -252 232 -76
rect -232 -580 -198 -404
rect -74 -580 -40 -404
rect 40 -580 74 -404
rect 198 -580 232 -404
<< poly >>
rect -186 673 -86 689
rect -186 639 -170 673
rect -102 639 -86 673
rect -186 592 -86 639
rect 86 673 186 689
rect 86 639 102 673
rect 170 639 186 673
rect 86 592 186 639
rect -186 345 -86 392
rect -186 311 -170 345
rect -102 311 -86 345
rect -186 264 -86 311
rect 86 345 186 392
rect 86 311 102 345
rect 170 311 186 345
rect 86 264 186 311
rect -186 17 -86 64
rect -186 -17 -170 17
rect -102 -17 -86 17
rect -186 -64 -86 -17
rect 86 17 186 64
rect 86 -17 102 17
rect 170 -17 186 17
rect 86 -64 186 -17
rect -186 -311 -86 -264
rect -186 -345 -170 -311
rect -102 -345 -86 -311
rect -186 -392 -86 -345
rect 86 -311 186 -264
rect 86 -345 102 -311
rect 170 -345 186 -311
rect 86 -392 186 -345
rect -186 -639 -86 -592
rect -186 -673 -170 -639
rect -102 -673 -86 -639
rect -186 -689 -86 -673
rect 86 -639 186 -592
rect 86 -673 102 -639
rect 170 -673 186 -639
rect 86 -689 186 -673
<< polycont >>
rect -170 639 -102 673
rect 102 639 170 673
rect -170 311 -102 345
rect 102 311 170 345
rect -170 -17 -102 17
rect 102 -17 170 17
rect -170 -345 -102 -311
rect 102 -345 170 -311
rect -170 -673 -102 -639
rect 102 -673 170 -639
<< locali >>
rect -186 639 -170 673
rect -102 639 -86 673
rect 86 639 102 673
rect 170 639 186 673
rect -232 580 -198 596
rect -232 388 -198 404
rect -74 580 -40 596
rect -74 388 -40 404
rect 40 580 74 596
rect 40 388 74 404
rect 198 580 232 596
rect 198 388 232 404
rect -186 311 -170 345
rect -102 311 -86 345
rect 86 311 102 345
rect 170 311 186 345
rect -232 252 -198 268
rect -232 60 -198 76
rect -74 252 -40 268
rect -74 60 -40 76
rect 40 252 74 268
rect 40 60 74 76
rect 198 252 232 268
rect 198 60 232 76
rect -186 -17 -170 17
rect -102 -17 -86 17
rect 86 -17 102 17
rect 170 -17 186 17
rect -232 -76 -198 -60
rect -232 -268 -198 -252
rect -74 -76 -40 -60
rect -74 -268 -40 -252
rect 40 -76 74 -60
rect 40 -268 74 -252
rect 198 -76 232 -60
rect 198 -268 232 -252
rect -186 -345 -170 -311
rect -102 -345 -86 -311
rect 86 -345 102 -311
rect 170 -345 186 -311
rect -232 -404 -198 -388
rect -232 -596 -198 -580
rect -74 -404 -40 -388
rect -74 -596 -40 -580
rect 40 -404 74 -388
rect 40 -596 74 -580
rect 198 -404 232 -388
rect 198 -596 232 -580
rect -186 -673 -170 -639
rect -102 -673 -86 -639
rect 86 -673 102 -639
rect 170 -673 186 -639
<< viali >>
rect -160 639 -112 673
rect 112 639 160 673
rect -232 404 -198 580
rect -74 404 -40 580
rect 40 404 74 580
rect 198 404 232 580
rect -160 311 -112 345
rect 112 311 160 345
rect -232 76 -198 252
rect -74 76 -40 252
rect 40 76 74 252
rect 198 76 232 252
rect -160 -17 -112 17
rect 112 -17 160 17
rect -232 -252 -198 -76
rect -74 -252 -40 -76
rect 40 -252 74 -76
rect 198 -252 232 -76
rect -160 -345 -112 -311
rect 112 -345 160 -311
rect -232 -580 -198 -404
rect -74 -580 -40 -404
rect 40 -580 74 -404
rect 198 -580 232 -404
rect -160 -673 -112 -639
rect 112 -673 160 -639
<< metal1 >>
rect -172 673 -100 679
rect -172 639 -160 673
rect -112 639 -100 673
rect -172 633 -100 639
rect 100 673 172 679
rect 100 639 112 673
rect 160 639 172 673
rect 100 633 172 639
rect -238 580 -192 592
rect -238 404 -232 580
rect -198 404 -192 580
rect -238 392 -192 404
rect -80 580 -34 592
rect -80 404 -74 580
rect -40 404 -34 580
rect -80 392 -34 404
rect 34 580 80 592
rect 34 404 40 580
rect 74 404 80 580
rect 34 392 80 404
rect 192 580 238 592
rect 192 404 198 580
rect 232 404 238 580
rect 192 392 238 404
rect -172 345 -100 351
rect -172 311 -160 345
rect -112 311 -100 345
rect -172 305 -100 311
rect 100 345 172 351
rect 100 311 112 345
rect 160 311 172 345
rect 100 305 172 311
rect -238 252 -192 264
rect -238 76 -232 252
rect -198 76 -192 252
rect -238 64 -192 76
rect -80 252 -34 264
rect -80 76 -74 252
rect -40 76 -34 252
rect -80 64 -34 76
rect 34 252 80 264
rect 34 76 40 252
rect 74 76 80 252
rect 34 64 80 76
rect 192 252 238 264
rect 192 76 198 252
rect 232 76 238 252
rect 192 64 238 76
rect -172 17 -100 23
rect -172 -17 -160 17
rect -112 -17 -100 17
rect -172 -23 -100 -17
rect 100 17 172 23
rect 100 -17 112 17
rect 160 -17 172 17
rect 100 -23 172 -17
rect -238 -76 -192 -64
rect -238 -252 -232 -76
rect -198 -252 -192 -76
rect -238 -264 -192 -252
rect -80 -76 -34 -64
rect -80 -252 -74 -76
rect -40 -252 -34 -76
rect -80 -264 -34 -252
rect 34 -76 80 -64
rect 34 -252 40 -76
rect 74 -252 80 -76
rect 34 -264 80 -252
rect 192 -76 238 -64
rect 192 -252 198 -76
rect 232 -252 238 -76
rect 192 -264 238 -252
rect -172 -311 -100 -305
rect -172 -345 -160 -311
rect -112 -345 -100 -311
rect -172 -351 -100 -345
rect 100 -311 172 -305
rect 100 -345 112 -311
rect 160 -345 172 -311
rect 100 -351 172 -345
rect -238 -404 -192 -392
rect -238 -580 -232 -404
rect -198 -580 -192 -404
rect -238 -592 -192 -580
rect -80 -404 -34 -392
rect -80 -580 -74 -404
rect -40 -580 -34 -404
rect -80 -592 -34 -580
rect 34 -404 80 -392
rect 34 -580 40 -404
rect 74 -580 80 -404
rect 34 -592 80 -580
rect 192 -404 238 -392
rect 192 -580 198 -404
rect 232 -580 238 -404
rect 192 -592 238 -580
rect -172 -639 -100 -633
rect -172 -673 -160 -639
rect -112 -673 -100 -639
rect -172 -679 -100 -673
rect 100 -639 172 -633
rect 100 -673 112 -639
rect 160 -673 172 -639
rect 100 -679 172 -673
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.5 m 4 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 70 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
