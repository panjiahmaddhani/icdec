magic
tech sky130A
magscale 1 2
timestamp 1729219847
<< nmos >>
rect -286 55 -86 455
rect 86 55 286 455
rect -286 -455 -86 -55
rect 86 -455 286 -55
<< ndiff >>
rect -344 443 -286 455
rect -344 67 -332 443
rect -298 67 -286 443
rect -344 55 -286 67
rect -86 443 -28 455
rect -86 67 -74 443
rect -40 67 -28 443
rect -86 55 -28 67
rect 28 443 86 455
rect 28 67 40 443
rect 74 67 86 443
rect 28 55 86 67
rect 286 443 344 455
rect 286 67 298 443
rect 332 67 344 443
rect 286 55 344 67
rect -344 -67 -286 -55
rect -344 -443 -332 -67
rect -298 -443 -286 -67
rect -344 -455 -286 -443
rect -86 -67 -28 -55
rect -86 -443 -74 -67
rect -40 -443 -28 -67
rect -86 -455 -28 -443
rect 28 -67 86 -55
rect 28 -443 40 -67
rect 74 -443 86 -67
rect 28 -455 86 -443
rect 286 -67 344 -55
rect 286 -443 298 -67
rect 332 -443 344 -67
rect 286 -455 344 -443
<< ndiffc >>
rect -332 67 -298 443
rect -74 67 -40 443
rect 40 67 74 443
rect 298 67 332 443
rect -332 -443 -298 -67
rect -74 -443 -40 -67
rect 40 -443 74 -67
rect 298 -443 332 -67
<< poly >>
rect -286 527 -86 543
rect -286 493 -270 527
rect -102 493 -86 527
rect -286 455 -86 493
rect 86 527 286 543
rect 86 493 102 527
rect 270 493 286 527
rect 86 455 286 493
rect -286 17 -86 55
rect -286 -17 -270 17
rect -102 -17 -86 17
rect -286 -55 -86 -17
rect 86 17 286 55
rect 86 -17 102 17
rect 270 -17 286 17
rect 86 -55 286 -17
rect -286 -493 -86 -455
rect -286 -527 -270 -493
rect -102 -527 -86 -493
rect -286 -543 -86 -527
rect 86 -493 286 -455
rect 86 -527 102 -493
rect 270 -527 286 -493
rect 86 -543 286 -527
<< polycont >>
rect -270 493 -102 527
rect 102 493 270 527
rect -270 -17 -102 17
rect 102 -17 270 17
rect -270 -527 -102 -493
rect 102 -527 270 -493
<< locali >>
rect -286 493 -270 527
rect -102 493 -86 527
rect 86 493 102 527
rect 270 493 286 527
rect -332 443 -298 459
rect -332 51 -298 67
rect -74 443 -40 459
rect -74 51 -40 67
rect 40 443 74 459
rect 40 51 74 67
rect 298 443 332 459
rect 298 51 332 67
rect -286 -17 -270 17
rect -102 -17 -86 17
rect 86 -17 102 17
rect 270 -17 286 17
rect -332 -67 -298 -51
rect -332 -459 -298 -443
rect -74 -67 -40 -51
rect -74 -459 -40 -443
rect 40 -67 74 -51
rect 40 -459 74 -443
rect 298 -67 332 -51
rect 298 -459 332 -443
rect -286 -527 -270 -493
rect -102 -527 -86 -493
rect 86 -527 102 -493
rect 270 -527 286 -493
<< viali >>
rect -245 493 -127 527
rect 127 493 245 527
rect -332 67 -298 443
rect -74 67 -40 443
rect 40 67 74 443
rect 298 67 332 443
rect -245 -17 -127 17
rect 127 -17 245 17
rect -332 -443 -298 -67
rect -74 -443 -40 -67
rect 40 -443 74 -67
rect 298 -443 332 -67
rect -245 -527 -127 -493
rect 127 -527 245 -493
<< metal1 >>
rect -257 527 -115 533
rect -257 493 -245 527
rect -127 493 -115 527
rect -257 487 -115 493
rect 115 527 257 533
rect 115 493 127 527
rect 245 493 257 527
rect 115 487 257 493
rect -338 443 -292 455
rect -338 67 -332 443
rect -298 67 -292 443
rect -338 55 -292 67
rect -80 443 -34 455
rect -80 67 -74 443
rect -40 67 -34 443
rect -80 55 -34 67
rect 34 443 80 455
rect 34 67 40 443
rect 74 67 80 443
rect 34 55 80 67
rect 292 443 338 455
rect 292 67 298 443
rect 332 67 338 443
rect 292 55 338 67
rect -257 17 -115 23
rect -257 -17 -245 17
rect -127 -17 -115 17
rect -257 -23 -115 -17
rect 115 17 257 23
rect 115 -17 127 17
rect 245 -17 257 17
rect 115 -23 257 -17
rect -338 -67 -292 -55
rect -338 -443 -332 -67
rect -298 -443 -292 -67
rect -338 -455 -292 -443
rect -80 -67 -34 -55
rect -80 -443 -74 -67
rect -40 -443 -34 -67
rect -80 -455 -34 -443
rect 34 -67 80 -55
rect 34 -443 40 -67
rect 74 -443 80 -67
rect 34 -455 80 -443
rect 292 -67 338 -55
rect 292 -443 298 -67
rect 332 -443 338 -67
rect 292 -455 338 -443
rect -257 -493 -115 -487
rect -257 -527 -245 -493
rect -127 -527 -115 -493
rect -257 -533 -115 -527
rect 115 -493 257 -487
rect 115 -527 127 -493
rect 245 -527 257 -493
rect 115 -533 257 -527
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 1 m 2 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 70 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
