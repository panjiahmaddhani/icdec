magic
tech sky130A
magscale 1 2
timestamp 1729241244
<< nwell >>
rect -552 -200 552 200
<< pmos >>
rect -458 -100 -358 100
rect -186 -100 -86 100
rect 86 -100 186 100
rect 358 -100 458 100
<< pdiff >>
rect -516 88 -458 100
rect -516 -88 -504 88
rect -470 -88 -458 88
rect -516 -100 -458 -88
rect -358 88 -300 100
rect -358 -88 -346 88
rect -312 -88 -300 88
rect -358 -100 -300 -88
rect -244 88 -186 100
rect -244 -88 -232 88
rect -198 -88 -186 88
rect -244 -100 -186 -88
rect -86 88 -28 100
rect -86 -88 -74 88
rect -40 -88 -28 88
rect -86 -100 -28 -88
rect 28 88 86 100
rect 28 -88 40 88
rect 74 -88 86 88
rect 28 -100 86 -88
rect 186 88 244 100
rect 186 -88 198 88
rect 232 -88 244 88
rect 186 -100 244 -88
rect 300 88 358 100
rect 300 -88 312 88
rect 346 -88 358 88
rect 300 -100 358 -88
rect 458 88 516 100
rect 458 -88 470 88
rect 504 -88 516 88
rect 458 -100 516 -88
<< pdiffc >>
rect -504 -88 -470 88
rect -346 -88 -312 88
rect -232 -88 -198 88
rect -74 -88 -40 88
rect 40 -88 74 88
rect 198 -88 232 88
rect 312 -88 346 88
rect 470 -88 504 88
<< poly >>
rect -458 181 -358 197
rect -458 147 -442 181
rect -374 147 -358 181
rect -458 100 -358 147
rect -186 181 -86 197
rect -186 147 -170 181
rect -102 147 -86 181
rect -186 100 -86 147
rect 86 181 186 197
rect 86 147 102 181
rect 170 147 186 181
rect 86 100 186 147
rect 358 181 458 197
rect 358 147 374 181
rect 442 147 458 181
rect 358 100 458 147
rect -458 -147 -358 -100
rect -458 -181 -442 -147
rect -374 -181 -358 -147
rect -458 -197 -358 -181
rect -186 -147 -86 -100
rect -186 -181 -170 -147
rect -102 -181 -86 -147
rect -186 -197 -86 -181
rect 86 -147 186 -100
rect 86 -181 102 -147
rect 170 -181 186 -147
rect 86 -197 186 -181
rect 358 -147 458 -100
rect 358 -181 374 -147
rect 442 -181 458 -147
rect 358 -197 458 -181
<< polycont >>
rect -442 147 -374 181
rect -170 147 -102 181
rect 102 147 170 181
rect 374 147 442 181
rect -442 -181 -374 -147
rect -170 -181 -102 -147
rect 102 -181 170 -147
rect 374 -181 442 -147
<< locali >>
rect -458 147 -442 181
rect -374 147 -358 181
rect -186 147 -170 181
rect -102 147 -86 181
rect 86 147 102 181
rect 170 147 186 181
rect 358 147 374 181
rect 442 147 458 181
rect -504 88 -470 104
rect -504 -104 -470 -88
rect -346 88 -312 104
rect -346 -104 -312 -88
rect -232 88 -198 104
rect -232 -104 -198 -88
rect -74 88 -40 104
rect -74 -104 -40 -88
rect 40 88 74 104
rect 40 -104 74 -88
rect 198 88 232 104
rect 198 -104 232 -88
rect 312 88 346 104
rect 312 -104 346 -88
rect 470 88 504 104
rect 470 -104 504 -88
rect -458 -181 -442 -147
rect -374 -181 -358 -147
rect -186 -181 -170 -147
rect -102 -181 -86 -147
rect 86 -181 102 -147
rect 170 -181 186 -147
rect 358 -181 374 -147
rect 442 -181 458 -147
<< viali >>
rect -442 147 -374 181
rect -170 147 -102 181
rect 102 147 170 181
rect 374 147 442 181
rect -504 -88 -470 88
rect -346 -88 -312 88
rect -232 -88 -198 88
rect -74 -88 -40 88
rect 40 -88 74 88
rect 198 -88 232 88
rect 312 -88 346 88
rect 470 -88 504 88
rect -442 -181 -374 -147
rect -170 -181 -102 -147
rect 102 -181 170 -147
rect 374 -181 442 -147
<< metal1 >>
rect -454 181 -362 187
rect -454 147 -442 181
rect -374 147 -362 181
rect -454 141 -362 147
rect -182 181 -90 187
rect -182 147 -170 181
rect -102 147 -90 181
rect -182 141 -90 147
rect 90 181 182 187
rect 90 147 102 181
rect 170 147 182 181
rect 90 141 182 147
rect 362 181 454 187
rect 362 147 374 181
rect 442 147 454 181
rect 362 141 454 147
rect -510 88 -464 100
rect -510 -88 -504 88
rect -470 -88 -464 88
rect -510 -100 -464 -88
rect -352 88 -306 100
rect -352 -88 -346 88
rect -312 -88 -306 88
rect -352 -100 -306 -88
rect -238 88 -192 100
rect -238 -88 -232 88
rect -198 -88 -192 88
rect -238 -100 -192 -88
rect -80 88 -34 100
rect -80 -88 -74 88
rect -40 -88 -34 88
rect -80 -100 -34 -88
rect 34 88 80 100
rect 34 -88 40 88
rect 74 -88 80 88
rect 34 -100 80 -88
rect 192 88 238 100
rect 192 -88 198 88
rect 232 -88 238 88
rect 192 -100 238 -88
rect 306 88 352 100
rect 306 -88 312 88
rect 346 -88 352 88
rect 306 -100 352 -88
rect 464 88 510 100
rect 464 -88 470 88
rect 504 -88 510 88
rect 464 -100 510 -88
rect -454 -147 -362 -141
rect -454 -181 -442 -147
rect -374 -181 -362 -147
rect -454 -187 -362 -181
rect -182 -147 -90 -141
rect -182 -181 -170 -147
rect -102 -181 -90 -147
rect -182 -187 -90 -181
rect 90 -147 182 -141
rect 90 -181 102 -147
rect 170 -181 182 -147
rect 90 -187 182 -181
rect 362 -147 454 -141
rect 362 -181 374 -147
rect 442 -181 454 -147
rect 362 -187 454 -181
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.5 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
