magic
tech sky130A
timestamp 1729132889
<< nwell >>
rect -97 -52 97 52
<< pmos >>
rect -50 -21 50 21
<< pdiff >>
rect -79 15 -50 21
rect -79 -15 -73 15
rect -56 -15 -50 15
rect -79 -21 -50 -15
rect 50 15 79 21
rect 50 -15 56 15
rect 73 -15 79 15
rect 50 -21 79 -15
<< pdiffc >>
rect -73 -15 -56 15
rect 56 -15 73 15
<< poly >>
rect -50 21 50 34
rect -50 -34 50 -21
<< locali >>
rect -73 15 -56 23
rect -73 -23 -56 -15
rect 56 15 73 23
rect 56 -23 73 -15
<< viali >>
rect -73 -15 -56 15
rect 56 -15 73 15
<< metal1 >>
rect -76 15 -53 21
rect -76 -15 -73 15
rect -56 -15 -53 15
rect -76 -21 -53 -15
rect 53 15 76 21
rect 53 -15 56 15
rect 73 -15 76 15
rect 53 -21 76 -15
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.42 l 1 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
